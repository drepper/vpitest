one.v