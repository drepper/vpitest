two.v